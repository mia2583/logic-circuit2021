-- Copyright (C) 2020  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and any partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details, at
-- https://fpgasoftware.intel.com/eula.

-- Generated by Quartus Prime Version 20.1.1 Build 720 11/11/2020 SJ Lite Edition
-- Created on Fri Nov 05 14:36:20 2021

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY CU IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        Din : IN STD_LOGIC_VECTOR(3 DOWNTO 0) := "0000";
        Dout : OUT STD_LOGIC
    );
END CU;

ARCHITECTURE BEHAVIOR OF CU IS
    TYPE type_fstate IS (state1,state2,state3,state4,state5);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,Din)
    BEGIN
        IF (reset='0') THEN
            reg_fstate <= state1;
            Dout <= '0';
        ELSE
            Dout <= '0';
            CASE fstate IS
                WHEN state1 =>
                    IF ((Din(3 DOWNTO 0) = "0011")) THEN
                        reg_fstate <= state2;
                    ELSIF ((Din(3 DOWNTO 0) /= "0011")) THEN
                        reg_fstate <= state1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state1;
                    END IF;

                    Dout <= '0';
                WHEN state2 =>
                    IF ((Din(3 DOWNTO 0) /= "1000")) THEN
                        reg_fstate <= state1;
                    ELSIF ((Din(3 DOWNTO 0) = "1000")) THEN
                        reg_fstate <= state3;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state2;
                    END IF;

                    Dout <= '0';
                WHEN state3 =>
                    IF ((Din(3 DOWNTO 0) /= "1001")) THEN
                        reg_fstate <= state1;
                    ELSIF ((Din(3 DOWNTO 0) = "1001")) THEN
                        reg_fstate <= state4;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state3;
                    END IF;

                    Dout <= '0';
                WHEN state4 =>
                    IF ((Din(3 DOWNTO 0) /= "0010")) THEN
                        reg_fstate <= state1;
                    ELSIF ((Din(3 DOWNTO 0) = "0010")) THEN
                        reg_fstate <= state5;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state4;
                    END IF;

                    Dout <= '0';
                WHEN state5 =>
                    IF ((Din(3 DOWNTO 0) /= "0011")) THEN
                        reg_fstate <= state1;
                    ELSIF ((Din(3 DOWNTO 0) = "0011")) THEN
                        reg_fstate <= state2;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state5;
                    END IF;

                    Dout <= '1';
                WHEN OTHERS => 
                    Dout <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
