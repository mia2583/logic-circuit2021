// Copyright (C) 2020  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// Generated by Quartus Prime Version 20.1.1 Build 720 11/11/2020 SJ Lite Edition
// Created on Wed Dec 22 16:10:43 2021

// synthesis message_off 10175

`timescale 1ns/1ns

module stop (
    reset,clock,same,way,
    nextFloor);

    input reset;
    input clock;
    input same;
    input way;

    output [3:0] nextFloor;
    reg [3:0] nextFloor;
    reg [8:0] fstate;
    reg [8:0] reg_fstate;
    parameter state1=0,state2=1,state3=2,state4=3,state6=4,state7=5,state8=6,state9=7,state5=8;

    always @(posedge clock)
    begin
        if (clock) begin
            fstate <= reg_fstate;
        end
    end

    always @(fstate or reset or same or way)
    begin
        if (~reset) begin
            reg_fstate <= state1;
            nextFloor <= 4'b0000;
        end
        else begin
            nextFloor <= 4'b0000;
            case (fstate)
                state1: begin
                    if (((way == 1'b1) & (same == 1'b0)))
                        reg_fstate <= state2;
                    else if ((way == 1'b0))
                        reg_fstate <= state1;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state1;

                    nextFloor <= 4'b0001;
                end
                state2: begin
                    if (((way == 1'b1) & (same == 1'b0)))
                        reg_fstate <= state3;
                    else if (((way == 1'b0) & (same == 1'b0)))
                        reg_fstate <= state1;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state2;

                    nextFloor <= 4'b0010;
                end
                state3: begin
                    if (((way == 1'b1) & (same == 1'b0)))
                        reg_fstate <= state4;
                    else if (((way == 1'b0) & (same == 1'b0)))
                        reg_fstate <= state2;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state3;

                    nextFloor <= 4'b0011;
                end
                state4: begin
                    if (((way == 1'b0) & (same == 1'b0)))
                        reg_fstate <= state3;
                    else if (((way == 1'b1) & (same == 1'b0)))
                        reg_fstate <= state5;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state4;

                    nextFloor <= 4'b0100;
                end
                state6: begin
                    if (((way == 1'b1) & (same == 1'b0)))
                        reg_fstate <= state7;
                    else if (((way == 1'b0) & (same == 1'b0)))
                        reg_fstate <= state5;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state6;

                    nextFloor <= 4'b0110;
                end
                state7: begin
                    if (((way == 1'b0) & (same == 1'b0)))
                        reg_fstate <= state6;
                    else if (((way == 1'b1) & (same == 1'b0)))
                        reg_fstate <= state8;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state7;

                    nextFloor <= 4'b0111;
                end
                state8: begin
                    if (((way == 1'b0) & (same == 1'b0)))
                        reg_fstate <= state7;
                    else if (((way == 1'b1) & (same == 1'b0)))
                        reg_fstate <= state9;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state8;

                    nextFloor <= 4'b1000;
                end
                state9: begin
                    if ((way == 1'b1))
                        reg_fstate <= state9;
                    else if (((way == 1'b0) & (same == 1'b0)))
                        reg_fstate <= state8;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state9;

                    nextFloor <= 4'b1001;
                end
                state5: begin
                    if (((way == 1'b0) & (same == 1'b0)))
                        reg_fstate <= state4;
                    else if (((way == 1'b1) & (same == 1'b0)))
                        reg_fstate <= state6;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state5;

                    nextFloor <= 4'b0101;
                end
                default: begin
                    nextFloor <= 4'bxxxx;
                    $display ("Reach undefined state");
                end
            endcase
        end
    end
endmodule // stop
